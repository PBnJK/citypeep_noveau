pBAV       ��       @       �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             �@             @;        ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��                @@         ��               L
�	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          